* File: adder.pex.sp
* Created: Sun Nov 10 00:17:27 2024
* Program "Calibre xRC"
* Version "v2022.3_33.19"
* 
.include "adder.pex.sp.pex"
.subckt adder  COUT A1 A2 A3 A4 B1 B2 B3 B4 CIN GND VDD S1 S2 S3 S4
* 
* S4	S4
* S3	S3
* S2	S2
* S1	S1
* VDD	VDD
* GND	GND
* CIN	CIN
* B4	B4
* B3	B3
* B2	B2
* B1	B1
* A4	A4
* A3	A3
* A2	A2
* A1	A1
* COUT	COUT
mXFA1/Mn14 N_C1_XFA1/Mn14_d N_XFA1/COB_XFA1/Mn14_g N_GND_XFA1/Mn14_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=1.4e-12 AS=1.5e-12 PD=3.8e-06
+ PS=4e-06
mXFA2/Mn14 N_C2_XFA2/Mn14_d N_XFA2/COB_XFA2/Mn14_g N_GND_XFA2/Mn14_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=1.4e-12 AS=1.5e-12 PD=3.8e-06
+ PS=4e-06
mXFA3/Mn14 N_C3_XFA3/Mn14_d N_XFA3/COB_XFA3/Mn14_g N_GND_XFA3/Mn14_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=1.4e-12 AS=1.5e-12 PD=3.8e-06
+ PS=4e-06
mXFA4/Mn14 N_COUT_XFA4/Mn14_d N_XFA4/COB_XFA4/Mn14_g N_GND_XFA4/Mn14_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=1.4e-12 AS=1.5e-12 PD=3.8e-06
+ PS=4e-06
mXFA1/Mn1 N_XFA1/N7_XFA1/Mn1_d N_A1_XFA1/Mn1_g N_GND_XFA1/Mn1_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=1.8e-12 AS=7e-13 PD=4.6e-06
+ PS=1.4e-06
mXFA2/Mn1 N_XFA2/N7_XFA2/Mn1_d N_A2_XFA2/Mn1_g N_GND_XFA2/Mn1_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=1.8e-12 AS=7e-13 PD=4.6e-06
+ PS=1.4e-06
mXFA3/Mn1 N_XFA3/N7_XFA3/Mn1_d N_A3_XFA3/Mn1_g N_GND_XFA3/Mn1_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=1.8e-12 AS=7e-13 PD=4.6e-06
+ PS=1.4e-06
mXFA4/Mn1 N_XFA4/N7_XFA4/Mn1_d N_A4_XFA4/Mn1_g N_GND_XFA4/Mn1_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=1.8e-12 AS=7e-13 PD=4.6e-06
+ PS=1.4e-06
mXFA1/Mn2 N_XFA1/N7_XFA1/Mn2_d N_B1_XFA1/Mn2_g N_GND_XFA1/Mn2_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA2/Mn2 N_XFA2/N7_XFA2/Mn2_d N_B2_XFA2/Mn2_g N_GND_XFA2/Mn2_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA3/Mn2 N_XFA3/N7_XFA3/Mn2_d N_B3_XFA3/Mn2_g N_GND_XFA3/Mn2_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA4/Mn2 N_XFA4/N7_XFA4/Mn2_d N_B4_XFA4/Mn2_g N_GND_XFA4/Mn2_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA1/Mn3 N_XFA1/COB_XFA1/Mn3_d N_CIN_XFA1/Mn3_g N_XFA1/N7_XFA1/Mn3_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA2/Mn3 N_XFA2/COB_XFA2/Mn3_d N_C1_XFA2/Mn3_g N_XFA2/N7_XFA2/Mn3_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA3/Mn3 N_XFA3/COB_XFA3/Mn3_d N_C2_XFA3/Mn3_g N_XFA3/N7_XFA3/Mn3_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA4/Mn3 N_XFA4/COB_XFA4/Mn3_d N_C3_XFA4/Mn3_g N_XFA4/N7_XFA4/Mn3_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA1/Mn5 N_XFA1/COB_XFA1/Mn5_d N_B1_XFA1/Mn5_g N_XFA1/N8_XFA1/Mn5_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA2/Mn5 N_XFA2/COB_XFA2/Mn5_d N_B2_XFA2/Mn5_g N_XFA2/N8_XFA2/Mn5_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA3/Mn5 N_XFA3/COB_XFA3/Mn5_d N_B3_XFA3/Mn5_g N_XFA3/N8_XFA3/Mn5_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA4/Mn5 N_XFA4/COB_XFA4/Mn5_d N_B4_XFA4/Mn5_g N_XFA4/N8_XFA4/Mn5_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA1/Mn4 N_XFA1/N8_XFA1/Mn4_d N_A1_XFA1/Mn4_g N_GND_XFA1/Mn4_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA2/Mn4 N_XFA2/N8_XFA2/Mn4_d N_A2_XFA2/Mn4_g N_GND_XFA2/Mn4_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA3/Mn4 N_XFA3/N8_XFA3/Mn4_d N_A3_XFA3/Mn4_g N_GND_XFA3/Mn4_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA4/Mn4 N_XFA4/N8_XFA4/Mn4_d N_A4_XFA4/Mn4_g N_GND_XFA4/Mn4_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA1/Mn6 N_XFA1/N9_XFA1/Mn6_d N_A1_XFA1/Mn6_g N_GND_XFA1/Mn6_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA2/Mn6 N_XFA2/N9_XFA2/Mn6_d N_A2_XFA2/Mn6_g N_GND_XFA2/Mn6_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA3/Mn6 N_XFA3/N9_XFA3/Mn6_d N_A3_XFA3/Mn6_g N_GND_XFA3/Mn6_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA4/Mn6 N_XFA4/N9_XFA4/Mn6_d N_A4_XFA4/Mn6_g N_GND_XFA4/Mn6_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA1/Mn7 N_XFA1/N9_XFA1/Mn7_d N_B1_XFA1/Mn7_g N_GND_XFA1/Mn7_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA2/Mn7 N_XFA2/N9_XFA2/Mn7_d N_B2_XFA2/Mn7_g N_GND_XFA2/Mn7_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA3/Mn7 N_XFA3/N9_XFA3/Mn7_d N_B3_XFA3/Mn7_g N_GND_XFA3/Mn7_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA4/Mn7 N_XFA4/N9_XFA4/Mn7_d N_B4_XFA4/Mn7_g N_GND_XFA4/Mn7_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA1/Mn8 N_XFA1/N9_XFA1/Mn8_d N_CIN_XFA1/Mn8_g N_GND_XFA1/Mn8_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA2/Mn8 N_XFA2/N9_XFA2/Mn8_d N_C1_XFA2/Mn8_g N_GND_XFA2/Mn8_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA3/Mn8 N_XFA3/N9_XFA3/Mn8_d N_C2_XFA3/Mn8_g N_GND_XFA3/Mn8_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA4/Mn8 N_XFA4/N9_XFA4/Mn8_d N_C3_XFA4/Mn8_g N_GND_XFA4/Mn8_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA1/Mn9 N_XFA1/SB_XFA1/Mn9_d N_XFA1/COB_XFA1/Mn9_g N_XFA1/N9_XFA1/Mn9_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA2/Mn9 N_XFA2/SB_XFA2/Mn9_d N_XFA2/COB_XFA2/Mn9_g N_XFA2/N9_XFA2/Mn9_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA3/Mn9 N_XFA3/SB_XFA3/Mn9_d N_XFA3/COB_XFA3/Mn9_g N_XFA3/N9_XFA3/Mn9_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA4/Mn9 N_XFA4/SB_XFA4/Mn9_d N_XFA4/COB_XFA4/Mn9_g N_XFA4/N9_XFA4/Mn9_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA1/Mn12 N_XFA1/SB_XFA1/Mn12_d N_CIN_XFA1/Mn12_g N_XFA1/N11_XFA1/Mn12_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA2/Mn12 N_XFA2/SB_XFA2/Mn12_d N_C1_XFA2/Mn12_g N_XFA2/N11_XFA2/Mn12_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA3/Mn12 N_XFA3/SB_XFA3/Mn12_d N_C2_XFA3/Mn12_g N_XFA3/N11_XFA3/Mn12_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA4/Mn12 N_XFA4/SB_XFA4/Mn12_d N_C3_XFA4/Mn12_g N_XFA4/N11_XFA4/Mn12_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA1/Mn11 N_XFA1/N11_XFA1/Mn11_d N_B1_XFA1/Mn11_g N_XFA1/N10_XFA1/Mn11_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA2/Mn11 N_XFA2/N11_XFA2/Mn11_d N_B2_XFA2/Mn11_g N_XFA2/N10_XFA2/Mn11_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA3/Mn11 N_XFA3/N11_XFA3/Mn11_d N_B3_XFA3/Mn11_g N_XFA3/N10_XFA3/Mn11_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA4/Mn11 N_XFA4/N11_XFA4/Mn11_d N_B4_XFA4/Mn11_g N_XFA4/N10_XFA4/Mn11_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA1/Mn10 N_XFA1/N10_XFA1/Mn10_d N_A1_XFA1/Mn10_g N_GND_XFA1/Mn10_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA2/Mn10 N_XFA2/N10_XFA2/Mn10_d N_A2_XFA2/Mn10_g N_GND_XFA2/Mn10_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA3/Mn10 N_XFA3/N10_XFA3/Mn10_d N_A3_XFA3/Mn10_g N_GND_XFA3/Mn10_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA4/Mn10 N_XFA4/N10_XFA4/Mn10_d N_A4_XFA4/Mn10_g N_GND_XFA4/Mn10_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=7e-13 AS=7e-13 PD=1.4e-06 PS=1.4e-06
mXFA1/Mn13 N_S1_XFA1/Mn13_d N_XFA1/SB_XFA1/Mn13_g N_GND_XFA1/Mn13_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=1.6e-12 AS=7e-13 PD=4.2e-06
+ PS=1.4e-06
mXFA2/Mn13 N_S2_XFA2/Mn13_d N_XFA2/SB_XFA2/Mn13_g N_GND_XFA2/Mn13_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=1.6e-12 AS=7e-13 PD=4.2e-06
+ PS=1.4e-06
mXFA3/Mn13 N_S3_XFA3/Mn13_d N_XFA3/SB_XFA3/Mn13_g N_GND_XFA3/Mn13_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=1.6e-12 AS=7e-13 PD=4.2e-06
+ PS=1.4e-06
mXFA4/Mn13 N_S4_XFA4/Mn13_d N_XFA4/SB_XFA4/Mn13_g N_GND_XFA4/Mn13_s
+ N_GND_XFA1/Mn14_b N_18 L=6e-07 W=1e-06 AD=1.6e-12 AS=7e-13 PD=4.2e-06
+ PS=1.4e-06
mXFA1/Mp14 N_C1_XFA1/Mp14_d N_XFA1/COB_XFA1/Mp14_g N_VDD_XFA1/Mp14_s
+ N_VDD_XFA1/Mp14_b P_18 L=6e-07 W=3e-06 AD=4.2e-12 AS=4.5e-12 PD=5.8e-06
+ PS=6e-06
mXFA2/Mp14 N_C2_XFA2/Mp14_d N_XFA2/COB_XFA2/Mp14_g N_VDD_XFA2/Mp14_s
+ N_VDD_XFA2/Mp14_b P_18 L=6e-07 W=3e-06 AD=4.2e-12 AS=4.5e-12 PD=5.8e-06
+ PS=6e-06
mXFA3/Mp14 N_C3_XFA3/Mp14_d N_XFA3/COB_XFA3/Mp14_g N_VDD_XFA3/Mp14_s
+ N_VDD_XFA3/Mp14_b P_18 L=6e-07 W=3e-06 AD=4.2e-12 AS=4.5e-12 PD=5.8e-06
+ PS=6e-06
mXFA4/Mp14 N_COUT_XFA4/Mp14_d N_XFA4/COB_XFA4/Mp14_g N_VDD_XFA4/Mp14_s
+ N_VDD_XFA4/Mp14_b P_18 L=6e-07 W=3e-06 AD=4.2e-12 AS=4.5e-12 PD=5.8e-06
+ PS=6e-06
mXFA1/Mp1 N_XFA1/N1_XFA1/Mp1_d N_A1_XFA1/Mp1_g N_VDD_XFA1/Mp1_s
+ N_VDD_XFA1/Mp14_b P_18 L=6e-07 W=3e-06 AD=5.4e-12 AS=2.1e-12 PD=6.6e-06
+ PS=1.4e-06
mXFA2/Mp1 N_XFA2/N1_XFA2/Mp1_d N_A2_XFA2/Mp1_g N_VDD_XFA2/Mp1_s
+ N_VDD_XFA2/Mp14_b P_18 L=6e-07 W=3e-06 AD=5.4e-12 AS=2.1e-12 PD=6.6e-06
+ PS=1.4e-06
mXFA3/Mp1 N_XFA3/N1_XFA3/Mp1_d N_A3_XFA3/Mp1_g N_VDD_XFA3/Mp1_s
+ N_VDD_XFA3/Mp14_b P_18 L=6e-07 W=3e-06 AD=5.4e-12 AS=2.1e-12 PD=6.6e-06
+ PS=1.4e-06
mXFA4/Mp1 N_XFA4/N1_XFA4/Mp1_d N_A4_XFA4/Mp1_g N_VDD_XFA4/Mp1_s
+ N_VDD_XFA4/Mp14_b P_18 L=6e-07 W=3e-06 AD=5.4e-12 AS=2.1e-12 PD=6.6e-06
+ PS=1.4e-06
mXFA1/Mp2 N_XFA1/N1_XFA1/Mp2_d N_B1_XFA1/Mp2_g N_VDD_XFA1/Mp2_s
+ N_VDD_XFA1/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA2/Mp2 N_XFA2/N1_XFA2/Mp2_d N_B2_XFA2/Mp2_g N_VDD_XFA2/Mp2_s
+ N_VDD_XFA2/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA3/Mp2 N_XFA3/N1_XFA3/Mp2_d N_B3_XFA3/Mp2_g N_VDD_XFA3/Mp2_s
+ N_VDD_XFA3/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA4/Mp2 N_XFA4/N1_XFA4/Mp2_d N_B4_XFA4/Mp2_g N_VDD_XFA4/Mp2_s
+ N_VDD_XFA4/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA1/Mp3 N_XFA1/COB_XFA1/Mp3_d N_CIN_XFA1/Mp3_g N_XFA1/N1_XFA1/Mp3_s
+ N_VDD_XFA1/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA2/Mp3 N_XFA2/COB_XFA2/Mp3_d N_C1_XFA2/Mp3_g N_XFA2/N1_XFA2/Mp3_s
+ N_VDD_XFA2/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA3/Mp3 N_XFA3/COB_XFA3/Mp3_d N_C2_XFA3/Mp3_g N_XFA3/N1_XFA3/Mp3_s
+ N_VDD_XFA3/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA4/Mp3 N_XFA4/COB_XFA4/Mp3_d N_C3_XFA4/Mp3_g N_XFA4/N1_XFA4/Mp3_s
+ N_VDD_XFA4/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA1/Mp5 N_XFA1/COB_XFA1/Mp5_d N_B1_XFA1/Mp5_g N_XFA1/N2_XFA1/Mp5_s
+ N_VDD_XFA1/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA2/Mp5 N_XFA2/COB_XFA2/Mp5_d N_B2_XFA2/Mp5_g N_XFA2/N2_XFA2/Mp5_s
+ N_VDD_XFA2/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA3/Mp5 N_XFA3/COB_XFA3/Mp5_d N_B3_XFA3/Mp5_g N_XFA3/N2_XFA3/Mp5_s
+ N_VDD_XFA3/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA4/Mp5 N_XFA4/COB_XFA4/Mp5_d N_B4_XFA4/Mp5_g N_XFA4/N2_XFA4/Mp5_s
+ N_VDD_XFA4/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA1/Mp4 N_XFA1/N2_XFA1/Mp4_d N_A1_XFA1/Mp4_g N_VDD_XFA1/Mp4_s
+ N_VDD_XFA1/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA2/Mp4 N_XFA2/N2_XFA2/Mp4_d N_A2_XFA2/Mp4_g N_VDD_XFA2/Mp4_s
+ N_VDD_XFA2/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA3/Mp4 N_XFA3/N2_XFA3/Mp4_d N_A3_XFA3/Mp4_g N_VDD_XFA3/Mp4_s
+ N_VDD_XFA3/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA4/Mp4 N_XFA4/N2_XFA4/Mp4_d N_A4_XFA4/Mp4_g N_VDD_XFA4/Mp4_s
+ N_VDD_XFA4/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA1/Mp6 N_XFA1/N3_XFA1/Mp6_d N_A1_XFA1/Mp6_g N_VDD_XFA1/Mp6_s
+ N_VDD_XFA1/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA2/Mp6 N_XFA2/N3_XFA2/Mp6_d N_A2_XFA2/Mp6_g N_VDD_XFA2/Mp6_s
+ N_VDD_XFA2/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA3/Mp6 N_XFA3/N3_XFA3/Mp6_d N_A3_XFA3/Mp6_g N_VDD_XFA3/Mp6_s
+ N_VDD_XFA3/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA4/Mp6 N_XFA4/N3_XFA4/Mp6_d N_A4_XFA4/Mp6_g N_VDD_XFA4/Mp6_s
+ N_VDD_XFA4/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA1/Mp7 N_XFA1/N3_XFA1/Mp7_d N_B1_XFA1/Mp7_g N_VDD_XFA1/Mp7_s
+ N_VDD_XFA1/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA2/Mp7 N_XFA2/N3_XFA2/Mp7_d N_B2_XFA2/Mp7_g N_VDD_XFA2/Mp7_s
+ N_VDD_XFA2/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA3/Mp7 N_XFA3/N3_XFA3/Mp7_d N_B3_XFA3/Mp7_g N_VDD_XFA3/Mp7_s
+ N_VDD_XFA3/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA4/Mp7 N_XFA4/N3_XFA4/Mp7_d N_B4_XFA4/Mp7_g N_VDD_XFA4/Mp7_s
+ N_VDD_XFA4/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA1/Mp8 N_XFA1/N3_XFA1/Mp8_d N_CIN_XFA1/Mp8_g N_VDD_XFA1/Mp8_s
+ N_VDD_XFA1/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA2/Mp8 N_XFA2/N3_XFA2/Mp8_d N_C1_XFA2/Mp8_g N_VDD_XFA2/Mp8_s
+ N_VDD_XFA2/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA3/Mp8 N_XFA3/N3_XFA3/Mp8_d N_C2_XFA3/Mp8_g N_VDD_XFA3/Mp8_s
+ N_VDD_XFA3/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA4/Mp8 N_XFA4/N3_XFA4/Mp8_d N_C3_XFA4/Mp8_g N_VDD_XFA4/Mp8_s
+ N_VDD_XFA4/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA1/Mp9 N_XFA1/SB_XFA1/Mp9_d N_XFA1/COB_XFA1/Mp9_g N_XFA1/N3_XFA1/Mp9_s
+ N_VDD_XFA1/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA2/Mp9 N_XFA2/SB_XFA2/Mp9_d N_XFA2/COB_XFA2/Mp9_g N_XFA2/N3_XFA2/Mp9_s
+ N_VDD_XFA2/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA3/Mp9 N_XFA3/SB_XFA3/Mp9_d N_XFA3/COB_XFA3/Mp9_g N_XFA3/N3_XFA3/Mp9_s
+ N_VDD_XFA3/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA4/Mp9 N_XFA4/SB_XFA4/Mp9_d N_XFA4/COB_XFA4/Mp9_g N_XFA4/N3_XFA4/Mp9_s
+ N_VDD_XFA4/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA1/Mp12 N_XFA1/SB_XFA1/Mp12_d N_CIN_XFA1/Mp12_g N_XFA1/N6_XFA1/Mp12_s
+ N_VDD_XFA1/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA2/Mp12 N_XFA2/SB_XFA2/Mp12_d N_C1_XFA2/Mp12_g N_XFA2/N6_XFA2/Mp12_s
+ N_VDD_XFA2/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA3/Mp12 N_XFA3/SB_XFA3/Mp12_d N_C2_XFA3/Mp12_g N_XFA3/N6_XFA3/Mp12_s
+ N_VDD_XFA3/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA4/Mp12 N_XFA4/SB_XFA4/Mp12_d N_C3_XFA4/Mp12_g N_XFA4/N6_XFA4/Mp12_s
+ N_VDD_XFA4/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA1/Mp11 N_XFA1/N6_XFA1/Mp11_d N_B1_XFA1/Mp11_g N_XFA1/N5_XFA1/Mp11_s
+ N_VDD_XFA1/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA2/Mp11 N_XFA2/N6_XFA2/Mp11_d N_B2_XFA2/Mp11_g N_XFA2/N5_XFA2/Mp11_s
+ N_VDD_XFA2/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA3/Mp11 N_XFA3/N6_XFA3/Mp11_d N_B3_XFA3/Mp11_g N_XFA3/N5_XFA3/Mp11_s
+ N_VDD_XFA3/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA4/Mp11 N_XFA4/N6_XFA4/Mp11_d N_B4_XFA4/Mp11_g N_XFA4/N5_XFA4/Mp11_s
+ N_VDD_XFA4/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA1/Mp10 N_XFA1/N5_XFA1/Mp10_d N_A1_XFA1/Mp10_g N_VDD_XFA1/Mp10_s
+ N_VDD_XFA1/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA2/Mp10 N_XFA2/N5_XFA2/Mp10_d N_A2_XFA2/Mp10_g N_VDD_XFA2/Mp10_s
+ N_VDD_XFA2/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA3/Mp10 N_XFA3/N5_XFA3/Mp10_d N_A3_XFA3/Mp10_g N_VDD_XFA3/Mp10_s
+ N_VDD_XFA3/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA4/Mp10 N_XFA4/N5_XFA4/Mp10_d N_A4_XFA4/Mp10_g N_VDD_XFA4/Mp10_s
+ N_VDD_XFA4/Mp14_b P_18 L=6e-07 W=3e-06 AD=2.1e-12 AS=2.1e-12 PD=1.4e-06
+ PS=1.4e-06
mXFA1/Mp13 N_S1_XFA1/Mp13_d N_XFA1/SB_XFA1/Mp13_g N_VDD_XFA1/Mp13_s
+ N_VDD_XFA1/Mp14_b P_18 L=6e-07 W=3e-06 AD=4.8e-12 AS=2.1e-12 PD=6.2e-06
+ PS=1.4e-06
mXFA2/Mp13 N_S2_XFA2/Mp13_d N_XFA2/SB_XFA2/Mp13_g N_VDD_XFA2/Mp13_s
+ N_VDD_XFA2/Mp14_b P_18 L=6e-07 W=3e-06 AD=4.8e-12 AS=2.1e-12 PD=6.2e-06
+ PS=1.4e-06
mXFA3/Mp13 N_S3_XFA3/Mp13_d N_XFA3/SB_XFA3/Mp13_g N_VDD_XFA3/Mp13_s
+ N_VDD_XFA3/Mp14_b P_18 L=6e-07 W=3e-06 AD=4.8e-12 AS=2.1e-12 PD=6.2e-06
+ PS=1.4e-06
mXFA4/Mp13 N_S4_XFA4/Mp13_d N_XFA4/SB_XFA4/Mp13_g N_VDD_XFA4/Mp13_s
+ N_VDD_XFA4/Mp14_b P_18 L=6e-07 W=3e-06 AD=4.8e-12 AS=2.1e-12 PD=6.2e-06
+ PS=1.4e-06
*
.include "adder.pex.sp.ADDER.pxi"
*
.ends
*
*
